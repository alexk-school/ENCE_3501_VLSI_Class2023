*** SPICE deck for cell dac{sch} from library lab1_dac
*** Created on Tue Sep 26, 2023 11:38:18
*** Last revised on Tue Sep 26, 2023 18:50:21
*** Written on Tue Sep 26, 2023 18:50:25 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT lab1_dac__div FROM CELL div{sch}
.SUBCKT lab1_dac__div bot in out
Rresnwell@0 net@0 in 10k
Rresnwell@1 out net@0 10k
Rresnwell@2 out bot 10k

* Spice Code nodes in cell cell 'div{sch}'
.ENDS lab1_dac__div

.global gnd

*** TOP LEVEL CELL: dac{sch}
Rresnwell@4 net@12 gnd 10k
Xdiv@0 net@1 b4 out lab1_dac__div
Xdiv@1 net@2 b3 net@1 lab1_dac__div
Xdiv@2 net@3 b2 net@2 lab1_dac__div
Xdiv@3 net@11 b1 net@3 lab1_dac__div
Xdiv@4 net@12 b0 net@11 lab1_dac__div

* Spice Code nodes in cell cell 'dac{sch}'
v4 b4 0
v3 b3 0
v2 b2 0
v1 b1 b0
vin b0 0 DC 5
.op
.END
