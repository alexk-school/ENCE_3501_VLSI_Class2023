*** SPICE deck for cell sim_2{sch} from library lab4
*** Created on Sun Oct 15, 2023 20:20:46
*** Last revised on Wed Oct 18, 2023 12:27:45
*** Written on Wed Oct 18, 2023 12:27:57 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT lab4__inverter_1 FROM CELL inverter_1{sch}
.SUBCKT lab4__inverter_1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 out in gnd gnd NMOS L=1.8U W=1.8U
Mpmos@2 out in vdd vdd PMOS L=1.8U W=3.6U
.ENDS lab4__inverter_1

*** SUBCIRCUIT lab4__inverter_2 FROM CELL inverter_2{sch}
.SUBCKT lab4__inverter_2 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 out in gnd gnd NMOS L=1.8U W=7.2U
Mpmos@0 out in vdd vdd PMOS L=1.8U W=14.4U
.ENDS lab4__inverter_2

.global gnd vdd

*** TOP LEVEL CELL: sim_2{sch}
Ccap@1 gnd vout2 {x}
Ccap@2 gnd vout1 {x}
Xinverter@0 vin vout1 lab4__inverter_1
Xinverter@2 vin vout2 lab4__inverter_2

* Spice Code nodes in cell cell 'sim_2{sch}'
vdd vdd 0 DC 5
vin vin 0 pulse(0v 5v 5n 1n 1n 12n 25n)
.step param x list 100f 1p 10p 100p
.trans 0 25n 0 100p
.include C5_models.txt
.END
