*** SPICE deck for cell ChargePump{sch} from library lab6
*** Created on Fri Nov 03, 2023 11:29:43
*** Last revised on Tue Nov 07, 2023 11:06:55
*** Written on Tue Nov 07, 2023 15:08:54 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: ChargePump{sch}
Ccap@0 OSC net@18 100u
Ccap@1 OSC2 net@6 100u
Ccap@2 OSC net@9 100u
Ccap@3 gnd Y 100u
Mnmos@0 vdd vdd net@18 gnd N_50n L=0.6U W=6U
Mnmos@6 net@18 net@18 net@6 gnd N_50n L=0.6U W=6U
Mnmos@7 net@6 net@6 net@9 gnd N_50n L=0.6U W=6U
Mnmos@8 net@9 net@9 Y gnd N_50n L=0.6U W=6U
Rresnwell@0 Y gnd 2MEG

* Spice Code nodes in cell cell 'ChargePump{sch}'
.include cmosedu_models.txt
vdd vdd 0 DC 1
v1 OSC 0 PULSE(0 1 0 1u 1u 12.5m 25m 1Meg)
v2 OSC2 0 PULSE(0 1 12.5m 1u 1u 12.5m 25m 1Meg)
.ic V(Y) = 0
.tran 0 100 0 20m
.END
